
module result_screen (
					input	logic clk,
					input	logic resetN,
					input logic	[10:0] pixelX,
					input logic	[10:0] pixelY,
					input logic win,
					input logic [3:0]lose,
					
					output	logic	drawingRequest,
					output	logic	[7:0] RGBout
);



localparam int WIDTH = 65;
localparam int HEIGHT = 16;

logic [0:HEIGHT-1] [0:WIDTH-1] win_bitmap = {
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b11101110001111110011100111000011100111001111100111001110000000000},
{65'b11101110011111111011100111000011100111001111100111001110000000000},
{65'b11101110011100111011100111000011100111000111000111101110000000000},
{65'b11101110011100111011100111000011100111000111000111111110000000000},
{65'b01111100011100111011100111000011100111000111000111111110000000000},
{65'b01111100011100111011100111000011111111000111000111111110000000000},
{65'b00111000011100111011100111000011111111000111000111011110000000000},
{65'b00111000011100111011100111000011111111000111000111001110000000000},
{65'b00111000011111111011111111000001100110001111100111001110000000000},
{65'b00111000001111110001111110000001100110001111100111001110000000000},
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b00000000000000000000000000000000000000000000000000000000000000000}
};

logic [0:HEIGHT-1] [0:WIDTH-1] lose_bitmap = {
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b11101110001111110011100111000011100000001111110001111110011111111},
{65'b11101110011111111011100111000011100000011111111011111111011111111},
{65'b11101110011100111011100111000011100000011100111011100111011100000},
{65'b11101110011100111011100111000011100000011100111011100000011100000},
{65'b01111100011100111011100111000011100000011100111011111110011111100},
{65'b01111100011100111011100111000011100000011100111001111111011111100},
{65'b00111000011100111011100111000011100000011100111000000111011100000},
{65'b00111000011100111011100111000011100000011100111011100111011100000},
{65'b00111000011111111011111111000011111111011111111011111111011111111},
{65'b00111000001111110001111110000011111111001111110001111110011111111},
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b00000000000000000000000000000000000000000000000000000000000000000},
{65'b00000000000000000000000000000000000000000000000000000000000000000}
};


localparam logic [10:0] topLeftX = 192;
localparam logic [10:0] topLeftY = 208;

logic signed [11:0] diffY;
logic signed [11:0] diffX;

localparam int SCALE_BITS = 2;

assign diffY = (pixelY - topLeftY) >> SCALE_BITS;
assign diffX = (pixelX - topLeftX) >> SCALE_BITS;

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
	end else begin
		drawingRequest = 0;

		if(0 <= diffX && diffX < WIDTH && diffY < HEIGHT) begin
			if(win == 1'b1) begin
				drawingRequest = win_bitmap[diffY][diffX];
			end else if(lose==0) begin
				drawingRequest = lose_bitmap[diffY][diffX];
			end
		end

		RGBout = 8'hFF;
	end
end

endmodule
